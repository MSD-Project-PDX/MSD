module top;
  logic mc_q[$:15];

  initial begin
    $display("dinesh_kumar size = %d,....%p",mc_q.size(), mc_q);
  end

endmodule
